module main

fn main() {
	server_init()
}
